module PC(PC_in,PC_out,RESET);
	input	[31:0]	PC_in;
	output	[31:0]	PC_out;
	input		RESET;

endmodule

module tb_MIPSALU2();
	
endmodule
